//////////////////////////////////////////////////////////////////////
//                                                                  //
//  File name : test_lib.svh                                        //
//  Author    : G. Andres Mancera                                   //
//  License   : GNU Lesser General Public License                   //
//  Course    : System and Functional Verification Using UVM        //
//              UCSC Silicon Valley Extension                       //
//                                                                  //
//////////////////////////////////////////////////////////////////////
`ifndef TEST_LIB__SVH
`define TEST_LIB__SVH

`include "bringup_packet_test.sv"
`include "oversized_packet_test.sv"
`include "undersized_packet_test.sv"
`include "small_large_packet_test.sv"
`include "small_ipg_packet_test.sv"
`include "zero_ipg_packet_test.sv"

`endif  // TEST_LIB__SVH
